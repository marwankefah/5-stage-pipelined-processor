
-- THE BUFFER BETWEEN MEMORY AND WRITEBACK


-- TODO COMPLETE THE BUFFER
-- [FIRST ATTEMPT AT PUSHING TO REPO]